`ifndef _scmp_alu_h
`define _scmp_alu_h

`define 	SCMP_ALU_ADD	4'd0
`define 	SCMP_ALU_SR	4'd1
`define 	SCMP_ALU_RRL	4'd2
`define 	SCMP_ALU_OR	4'd3
`define 	SCMP_ALU_AND	4'd4
`define 	SCMP_ALU_XOR	4'd5
`define 	SCMP_ALU_INC	4'd6
`define 	SCMP_ALU_DEC	4'd7

`endif