`ifndef _scmp_microcode_h_
`define _scmp_microcode_h_

`include "scmp_microcode_pla.gen.vh"


`endif