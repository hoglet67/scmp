`ifndef _scmp_alu_h
`define _scmp_alu_h

`define 	SZ_ALU_OP	4
`define 	ALU_OP_ADD	4'd0
`define 	ALU_OP_SR	4'd1
`define 	ALU_OP_RRL	4'd2
`define 	ALU_OP_OR	4'd3
`define 	ALU_OP_AND	4'd4
`define 	ALU_OP_XOR	4'd5
`define 	ALU_OP_INC	4'd6
`define 	ALU_OP_DEC	4'd7
`define 	ALU_OP_NUL	`ALU_OP_INC

`endif